----------------------------------------------------------------------------------
-- Company: Esigelec
-- Engineer: Yash Motagi
-- 
-- Create Date:    06:39:01 06/12/2018 
-- Design Name: 
-- Module Name:    piccolokey - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity piccolokey is
generic( round : integer range 0 to 32
			);
port ( keyin : in std_logic_vector (127 downto 0);
		 key_out1_wk : out std_logic_vector (15 downto 0);
		 key_out2_wk : out std_logic_vector (15 downto 0);
		 key_out1_rk : out std_logic_vector (15 downto 0);
		 key_out2_rk : out std_logic_vector (15 downto 0));
end piccolokey;

architecture Behavioral of piccolokey is

component rk is
generic( round : integer range 0 to 32
			);
port ( key_in : in std_logic_vector (127 downto 0);
		 key_out_rk1 : out std_logic_vector (15 downto 0);
		 key_out_rk2 : out std_logic_vector (15 downto 0));
end component rk;

component wk is
generic( round : integer range 0 to 32
			);
port ( key_in : in std_logic_vector (127 downto 0);
		 key_out1_wk : out std_logic_vector (15 downto 0);
		 key_out2_wk : out std_logic_vector (15 downto 0));
end component wk;

component constant_gen is
generic( round : integer range 0 to 32
			);
port ( con : out std_logic_vector (31 downto 0));
end component constant_gen;

signal rk_1,rk_2 : std_logic_vector (15 downto 0);
signal const : std_logic_vector (31 downto 0);
begin

rk_component : rk
generic map( round => round
			)
port map( key_in => keyin,
		 key_out_rk1 =>rk_1,
		 key_out_rk2 =>rk_2);

wk_component : wk
generic map( round => round
			)
port map( key_in => keyin,
			 key_out1_wk => key_out1_wk,
			 key_out2_wk => key_out2_wk);
			 
constant_component : constant_gen
generic map( round => round
			)
port map( con => const);

out_process : process (keyin) is
begin
	key_out1_rk <= rk_1 xor const(31 downto 16);
	key_out2_rk <=	rk_2 xor const(15 downto 0);
end process	out_process;
	
end Behavioral;
